// PLL.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module PLL (
		input  wire  clkin_clk,   //   clkin.clk
		output wire  clkout1_clk, // clkout1.clk
		output wire  clkout2_clk, // clkout2.clk
		input  wire  reset_reset  //   reset.reset
	);

	PLL_altpll_0 altpll_0 (
		.clk       (clkin_clk),   //       inclk_interface.clk
		.reset     (reset_reset), // inclk_interface_reset.reset
		.read      (),            //             pll_slave.read
		.write     (),            //                      .write
		.address   (),            //                      .address
		.readdata  (),            //                      .readdata
		.writedata (),            //                      .writedata
		.c0        (clkout1_clk), //                    c0.clk
		.c1        (clkout2_clk)  //                    c1.clk
	);

endmodule
